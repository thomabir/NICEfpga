module CordicFSR #(
    parameter int BIT_WIDTH = 24
) (
    input logic clk_i,  // clock
    input logic start_i,  // start the computation
    input logic [BIT_WIDTH-1:0] sin_in,  // sine
    input logic [BIT_WIDTH-1:0] cos_in,  // cosine
    output logic [BIT_WIDTH-1:0] phi_out,  // phase
    output logic done_o  // computation is done, result is valid
);

    parameter int ITER = $clog2(BIT_WIDTH) + 1;  // 24 bit numbers -> 5 bit counter

    // CORDIC rotation angles in radians
    // Calculate the scale factor for angle values based on the number of iterations and bitwidth
    localparam ANGLE_SCALE = 1 << (BIT_WIDTH - 1);

    // Generate CORDIC rotation angles in radians at compile time
    genvar j;
    for (j = 0; j <= ITER; j = j + 1) begin
        localparam angle[i] = ANGLE_SCALE * $arctan(2 ** (-i));
    end


    typedef enum logic [2:0] {
        IDLE,  // wait for start_i, all outputs are zero
        ITERATE,  // iterate the CORDIC algorithm for BIT_WIDTH iterations
        DONE  // phi_out is valid, done_o is high, go back to IDLE
    } state_e;

    typedef struct packed {
        state_e state;
        logic [ITER-1:0] i;  // counts from BIT_WIDTH-1 to 0
        logic [BIT_WIDTH-1:0] x;  // x coordinate
        logic [BIT_WIDTH-1:0] y;  // y coordinate
        logic [BIT_WIDTH-1:0] phi;  // phase
        logic [BIT_WIDTH-1:0] phi_final;  // final phase, always valid
    } state_t;

    state_t state_d;
    state_t state_q;

    // start routine
    always_ff @(posedge clk_i) begin
        if (start_i) state_q.state <= IDLE;
        else state_q <= state_d;
    end  // always_ff


    always_comb begin
        state_d = state_q;

        case (state_q.state)

            // take inputs, get ready for computation
            IDLE: begin
                state_d.i = ITER'(BIT_WIDTH - 1);  // 23
                state_d.x = sin_in;
                state_d.y = cos_in;
                state_d.phi = 0;
                if (start_i) state_d.state = ITERATE;
            end

            ITERATE: begin
                if (state_q.i == 0) begin
                    state_d.state = DONE;
                    state_d.phi_final = state_q.phi;
                end
                else begin
                    if (state_q.x >= 0) begin
                        state_d.x = state_q.x - (state_q.y >>> state_q.i);
                        state_d.y = state_q.y + (state_q.x >>> state_q.i);
                        state_d.phi = state_q.phi + angle[state_q.i];
                    end
                    else begin
                        state_d.x = state_q.x + (state_q.y >>> state_q.i);
                        state_d.y = state_q.y - (state_q.x >>> state_q.i);
                        state_d.phi = state_q.phi - angle[state_q.i];
                    end
                    state_d.i = state_q.i - 1;
                end

            end

            DONE: begin
                state_d.state = IDLE;
            end

            default: begin
                state_d.state = IDLE;
            end

        endcase

        // output signals
        phi_out = state_q.phi_final;
        done_o = (state_q.state == DONE);


    end  // always_comb

endmodule
